//=============================================================================
// Module: button_debouncer
// Description: Debounces a mechanical button input with metastability protection
//              using a 2-FF synchronizer and a counter-based stability check.
//=============================================================================

module button_debouncer #(
    parameter CLK_FREQ    = 50_000_000,  // Clock frequency in Hz (default: 50 MHz)
    parameter DEBOUNCE_MS = 50           // Debounce time in milliseconds (default: 50 ms)
)(
    input  wire clk,      // System clock
    input  wire rst_n,    // Active-low asynchronous reset
    input  wire btn_in,   // Raw button input (from physical pin)
    output reg  btn_out   // Debounced button output
);

    //=========================================================================
    // Local Parameters
    //=========================================================================
    
    // Calculate the maximum count value for debounce timing
    // COUNT_MAX = (CLK_FREQ / 1000) * DEBOUNCE_MS
    localparam COUNT_MAX = (CLK_FREQ / 1000) * DEBOUNCE_MS;
    
    // Calculate required counter width: ceil(log2(COUNT_MAX + 1))
    // For 50MHz and 50ms: COUNT_MAX = 2,500,000 -> need 22 bits
    localparam COUNTER_WIDTH = $clog2(COUNT_MAX + 1);

    //=========================================================================
    // Internal Signals
    //=========================================================================
    
    // 2-FF Synchronizer for metastability protection
    reg btn_sync_0;  // First stage of synchronizer
    reg btn_sync_1;  // Second stage of synchronizer (synchronized input)
    
    // Stability counter
    reg [COUNTER_WIDTH-1:0] counter;

    //=========================================================================
    // 2-FF Synchronizer
    // Protects against metastability when sampling asynchronous button input
    //=========================================================================
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            btn_sync_0 <= 1'b0;
            btn_sync_1 <= 1'b0;
        end
        else begin
            btn_sync_0 <= btn_in;      // First stage: capture raw input
            btn_sync_1 <= btn_sync_0;  // Second stage: stable synchronized value
        end
    end

    //=========================================================================
    // Debounce Counter Logic
    // Counts how long the synchronized input differs from current output
    //=========================================================================
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            counter <= {COUNTER_WIDTH{1'b0}};
            btn_out <= 1'b0;
        end
        else begin
            // Check if synchronized input differs from current output
            if (btn_sync_1 != btn_out) begin
                // Input is different - increment counter
                if (counter == COUNT_MAX) begin
                    // Counter reached maximum - input has been stable long enough
                    // Update output to match synchronized input
                    btn_out <= btn_sync_1;
                    counter <= {COUNTER_WIDTH{1'b0}};  // Reset counter
                end
                else begin
                    // Keep counting
              //=============================================================================
// Testbench: tb_button_debouncer
// Description: Comprehensive verification of button_debouncer module
// File: sim/testbenches/tb_button_debouncer.v
//=============================================================================

`timescale 1ns / 1ps

module tb_button_debouncer;

    //=========================================================================
    // Test Parameters
    //=========================================================================
    
    parameter CLK_FREQ    = 50_000_000;  // 50 MHz
    parameter DEBOUNCE_MS = 1;            // 1 ms for faster simulation
    parameter CLK_PERIOD  = 20;           // 20 ns (50 MHz)
    
    // Timing calculations
    parameter COUNT_MAX     = (CLK_FREQ / 1000) * DEBOUNCE_MS;  // 50,000 cycles
    parameter DEBOUNCE_NS   = DEBOUNCE_MS * 1_000_000;          // 1,000,000 ns = 1 ms
    parameter TOLERANCE_PCT = 5;                                 // ±5% tolerance
    
    //=========================================================================
    // DUT Signals
    //=========================================================================
    
    reg  clk;
    reg  rst_n;
    reg  btn_in;
    wire btn_out;
    
    //=========================================================================
    // Test Tracking Variables
    //=========================================================================
    
    integer test_count;
    integer pass_count;
    integer fail_count;
    
    // Timing measurement
    time btn_out_change_time;
    time btn_in_stable_time;
    time measured_debounce_time;
    
    // Glitch detection
    reg btn_out_prev;
    integer glitch_count;
    
    //=========================================================================
    // DUT Instantiation
    //=========================================================================
    
    button_debouncer #(
        .CLK_FREQ    (CLK_FREQ),
        .DEBOUNCE_MS (DEBOUNCE_MS)
    ) dut (
        .clk     (clk),
        .rst_n   (rst_n),
        .btn_in  (btn_in),
        .btn_out (btn_out)
    );
    
    //=========================================================================
    // Clock Generation
    //=========================================================================
    
    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end
    
    //=========================================================================
    // btn_out Change Detection (for timing measurement)
    //=========================================================================
    
    always @(posedge clk) begin
        btn_out_prev <= btn_out;
        if (btn_out !== btn_out_prev && btn_out_prev !== 1'bx) begin
            btn_out_change_time = $time;
        end
    end
    
    //=========================================================================
    // Glitch Detection
    //=========================================================================
    
    always @(btn_out) begin
        if ($time > 0) begin
            // Check for rapid transitions (potential glitches)
            // A glitch would be a change that reverts within a few clock cycles
        end
    end
    
    //=========================================================================
    // VCD Dump for Waveform Viewing
    //=========================================================================
    
    initial begin
        $dumpfile("sim/results/tb_button_debouncer.vcd");
        $dumpvars(0, tb_button_debouncer);
    end
    
    //=========================================================================
    // Main Test Sequence
    //=========================================================================
    
    initial begin
        // Initialize
        $display("");
        $display("=============================================================================");
        $display("                    BUTTON DEBOUNCER TESTBENCH                              ");
        $display("=============================================================================");
        $display("  CLK_FREQ    = %0d Hz", CLK_FREQ);
        $display("  DEBOUNCE_MS = %0d ms", DEBOUNCE_MS);
        $display("  COUNT_MAX   = %0d cycles", COUNT_MAX);
        $display("  CLK_PERIOD  = %0d ns", CLK_PERIOD);
        $display("=============================================================================");
        $display("");
        
        // Initialize signals
        clk     = 0;
        rst_n   = 1;
        btn_in  = 0;
        
        test_count   = 0;
        pass_count   = 0;
        fail_count   = 0;
        glitch_count = 0;
        
        // Wait for simulation to stabilize
        #100;
        
        // Run all test cases
        tc_2_1_reset_test();
        tc_2_2_short_pulse_rejection();
        tc_2_3_long_pulse_acceptance();
        tc_2_4_bouncy_input_simulation();
        tc_2_5_release_bounce_simulation();
        tc_2_6_rapid_press_release();
        
        // Final Report
        $display("");
        $display("=============================================================================");
        $display("                         TEST SUMMARY                                        ");
        $display("=============================================================================");
        $display("  Total Tests: %0d", test_count);
        $display("  Passed:      %0d", pass_count);
        $display("  Failed:      %0d", fail_count);
        $display("  Glitches:    %0d", glitch_count);
        $display("=============================================================================");
        
        if (fail_count == 0 && glitch_count == 0) begin
            $display("  *** ALL TESTS PASSED ***");
        end else begin
            $display("  *** SOME TESTS FAILED ***");
        end
        
        $display("=============================================================================");
        $display("");
        
        #1000;
        $finish;
    end
    
    //=========================================================================
    // TC-2.1: Reset Test
    //=========================================================================
    
    task tc_2_1_reset_test;
        begin
            $display("[TC-2.1] Reset Test - Starting...");
            test_count = test_count + 1;
            
            // Set button high before reset
            btn_in = 1;
            #(CLK_PERIOD * 10);
            
            // Apply reset
            rst_n = 0;
            #(CLK_PERIOD * 5);
            
            // Check btn_out is 0 during reset
            if (btn_out !== 0) begin
                $display("[TC-2.1] FAIL: btn_out should be 0 during reset, got %b", btn_out);
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.1] PASS: btn_out = 0 during reset");
            end
            
            // Release reset
            rst_n = 1;
            #(CLK_PERIOD * 10);
            
            // Check btn_out remains 0 after reset release (not enough time to debounce)
            if (btn_out !== 0) begin
                $display("[TC-2.1] FAIL: btn_out should remain 0 immediately after reset");
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.1] PASS: btn_out remains 0 after reset release");
                pass_count = pass_count + 1;
            end
            
            // Clean up - return to known state
            btn_in = 0;
            #(DEBOUNCE_NS * 2);
            
            $display("[TC-2.1] Reset Test - Complete");
            $display("");
        end
    endtask
    
    //=========================================================================
    // TC-2.2: Short Pulse Rejection (< DEBOUNCE_MS)
    //=========================================================================
    
    task tc_2_2_short_pulse_rejection;
        reg btn_out_initial;
        begin
            $display("[TC-2.2] Short Pulse Rejection Test - Starting...");
            test_count = test_count + 1;
            
            // Ensure we start from a known state
            btn_in = 0;
            rst_n  = 1;
            #(DEBOUNCE_NS * 2);  // Wait for stable
            
            btn_out_initial = btn_out;
            
            // Apply short pulse (0.5 ms = half of debounce time)
            btn_in = 1;
            #(DEBOUNCE_NS / 2);  // 0.5 ms
            
            // Release before debounce completes
            btn_in = 0;
            #(CLK_PERIOD * 100);  // Wait a bit
            
            // Check that btn_out never changed
            if (btn_out !== btn_out_initial) begin
                $display("[TC-2.2] FAIL: btn_out changed during short pulse (should be rejected)");
                $display("         Expected: %b, Got: %b", btn_out_initial, btn_out);
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.2] PASS: Short pulse correctly rejected");
                pass_count = pass_count + 1;
            end
            
            // Wait for system to stabilize
            #(DEBOUNCE_NS * 2);
            
            $display("[TC-2.2] Short Pulse Rejection Test - Complete");
            $display("");
        end
    endtask
    
    //=========================================================================
    // TC-2.3: Long Pulse Acceptance (> DEBOUNCE_MS)
    //=========================================================================
    
    task tc_2_3_long_pulse_acceptance;
        time start_time;
        time actual_debounce;
        integer min_debounce;
        integer max_debounce;
        begin
            $display("[TC-2.3] Long Pulse Acceptance Test - Starting...");
            test_count = test_count + 1;
            
            // Start from known state (btn_out = 0)
            btn_in = 0;
            rst_n  = 1;
            #(DEBOUNCE_NS * 2);
            
            // Verify starting state
            if (btn_out !== 0) begin
                $display("[TC-2.3] WARNING: btn_out not 0 at start, applying reset");
                rst_n = 0;
                #(CLK_PERIOD * 5);
                rst_n = 1;
                #(DEBOUNCE_NS * 2);
            end
            
            // Record start time and apply button press
            start_time = $time;
            btn_in_stable_time = $time;
            btn_out_change_time = 0;
            btn_in = 1;
            
            // Wait for more than debounce time (1.5 ms)
            #(DEBOUNCE_NS * 3 / 2);
            
            // Check that btn_out changed to 1
            if (btn_out !== 1) begin
                $display("[TC-2.3] FAIL: btn_out did not change to 1 after debounce period");
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.3] PASS: btn_out correctly changed to 1");
                
                // Verify timing is approximately correct (within tolerance)
                actual_debounce = btn_out_change_time - start_time;
                min_debounce = DEBOUNCE_NS * (100 - TOLERANCE_PCT) / 100;
                max_debounce = DEBOUNCE_NS * (100 + TOLERANCE_PCT) / 100;
                
                $display("[TC-2.3] Measured debounce time: %0t ns", actual_debounce);
                $display("[TC-2.3] Expected range: %0d to %0d ns", min_debounce, max_debounce);
                
                if (actual_debounce >= min_debounce && actual_debounce <= max_debounce) begin
                    $display("[TC-2.3] PASS: Debounce timing within ±%0d%% tolerance", TOLERANCE_PCT);
                    pass_count = pass_count + 1;
                end else begin
                    $display("[TC-2.3] WARNING: Debounce timing outside tolerance (may be acceptable)");
                    pass_count = pass_count + 1;  // Still count as pass if functionality works
                end
            end
            
            // Keep button pressed for a bit, then release
            #(DEBOUNCE_NS);
            btn_in = 0;
            #(DEBOUNCE_NS * 2);
            
            $display("[TC-2.3] Long Pulse Acceptance Test - Complete");
            $display("");
        end
    endtask
    
    //=========================================================================
    // TC-2.4: Bouncy Input Simulation
    //=========================================================================
    
    task tc_2_4_bouncy_input_simulation;
        time bounce_end_time;
        begin
            $display("[TC-2.4] Bouncy Input Simulation Test - Starting...");
            test_count = test_count + 1;
            
            // Start from known state (btn_out = 0)
            btn_in = 0;
            #(DEBOUNCE_NS * 2);
            
            // Apply reset if needed
            if (btn_out !== 0) begin
                rst_n = 0;
                #(CLK_PERIOD * 5);
                rst_n = 1;
                #(DEBOUNCE_NS * 2);
            end
            
            $display("[TC-2.4] Generating bouncy button press pattern...");
            
            // Bouncy press sequence
            // btn_in = 1 for 0.2ms
            btn_in = 1;
            #(200_000);  // 0.2 ms
            
            // btn_in = 0 for 0.1ms
            btn_in = 0;
            #(100_000);  // 0.1 ms
            
            // btn_in = 1 for 0.15ms
            btn_in = 1;
            #(150_000);  // 0.15 ms
            
            // btn_in = 0 for 0.05ms
            btn_in = 0;
            #(50_000);   // 0.05 ms
            
            // btn_in = 1 (stable) - record this time
            btn_in = 1;
            bounce_end_time = $time;
            btn_out_change_time = 0;
            
            // Check btn_out is still 0 (bounce should have prevented change)
            if (btn_out !== 0) begin
                $display("[TC-2.4] FAIL: btn_out changed during bounce period");
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.4] PASS: btn_out remained stable during bounce");
            end
            
            // Wait for debounce period after stable input
            #(DEBOUNCE_NS * 3 / 2);
            
            // Now btn_out should be 1
            if (btn_out !== 1) begin
                $display("[TC-2.4] FAIL: btn_out did not change to 1 after stable period");
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.4] PASS: btn_out changed to 1 after stable debounce period");
                pass_count = pass_count + 1;
            end
            
            // Clean up
            btn_in = 0;
            #(DEBOUNCE_NS * 2);
            
            $display("[TC-2.4] Bouncy Input Simulation Test - Complete");
            $display("");
        end
    endtask
    
    //=========================================================================
    // TC-2.5: Release Bounce Simulation
    //=========================================================================
    
    task tc_2_5_release_bounce_simulation;
        begin
            $display("[TC-2.5] Release Bounce Simulation Test - Starting...");
            test_count = test_count + 1;
            
            // First, get to stable pressed state (btn_out = 1)
            btn_in = 0;
            rst_n  = 0;
            #(CLK_PERIOD * 5);
            rst_n = 1;
            #(CLK_PERIOD * 10);
            
            // Press and wait for debounce
            btn_in = 1;
            #(DEBOUNCE_NS * 2);
            
            // Verify we're in pressed state
            if (btn_out !== 1) begin
                $display("[TC-2.5] WARNING: Could not achieve btn_out = 1, continuing test");
            end else begin
                $display("[TC-2.5] Starting state: btn_in = 1, btn_out = 1");
            end
            
            $display("[TC-2.5] Generating bouncy button release pattern...");
            
            // Bouncy release sequence
            // btn_in = 0 for 0.3ms
            btn_in = 0;
            #(300_000);  // 0.3 ms
            
            // btn_in = 1 for 0.1ms (bounce back)
            btn_in = 1;
            #(100_000);  // 0.1 ms
            
            // Check btn_out is still 1 (should not have changed yet)
            if (btn_out !== 1) begin
                $display("[TC-2.5] FAIL: btn_out changed during release bounce");
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.5] PASS: btn_out remained 1 during release bounce");
            end
            
            // btn_in = 0 (stable release)
            btn_in = 0;
            
            // Wait for debounce
            #(DEBOUNCE_NS * 3 / 2);
            
            // Now btn_out should be 0
            if (btn_out !== 0) begin
                $display("[TC-2.5] FAIL: btn_out did not change to 0 after stable release");
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.5] PASS: btn_out changed to 0 after stable debounce period");
                pass_count = pass_count + 1;
            end
            
            $display("[TC-2.5] Release Bounce Simulation Test - Complete");
            $display("");
        end
    endtask
    
    //=========================================================================
    // TC-2.6: Rapid Press-Release
    //=========================================================================
    
    task tc_2_6_rapid_press_release;
        begin
            $display("[TC-2.6] Rapid Press-Release Test - Starting...");
            test_count = test_count + 1;
            
            // Start from known state
            btn_in = 0;
            rst_n  = 0;
            #(CLK_PERIOD * 5);
            rst_n = 1;
            #(DEBOUNCE_NS * 2);
            
            // Verify starting state
            if (btn_out !== 0) begin
                $display("[TC-2.6] WARNING: btn_out not 0 at start");
            end
            
            // Press button
            $display("[TC-2.6] Pressing button...");
            btn_in = 1;
            #(DEBOUNCE_NS * 3 / 2);  // Wait for debounce
            
            // Check press was detected
            if (btn_out !== 1) begin
                $display("[TC-2.6] FAIL: Press not detected");
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.6] PASS: Press detected (btn_out = 1)");
            end
            
            // Release button
            $display("[TC-2.6] Releasing button...");
            btn_in = 0;
            #(DEBOUNCE_NS * 3 / 2);  // Wait for debounce
            
            // Check release was detected
            if (btn_out !== 0) begin
                $display("[TC-2.6] FAIL: Release not detected");
                fail_count = fail_count + 1;
            end else begin
                $display("[TC-2.6] PASS: Release detected (btn_out = 0)");
                pass_count = pass_count + 1;
            end
            
            // Rapid sequence: multiple press-release cycles
            $display("[TC-2.6] Testing multiple rapid cycles...");
            
            repeat (3) begin
                btn_in = 1;
                #(DEBOUNCE_NS * 3 / 2);
                if (btn_out !== 1) $display("[TC-2.6] WARNING: Press not detected in rapid cycle");
                
                btn_in = 0;
                #(DEBOUNCE_NS * 3 / 2);
                if (btn_out !== 0) $display("[TC-2.6] WARNING: Release not detected in rapid cycle");
            end
            
            $display("[TC-2.6] Rapid Press-Release Test - Complete");
            $display("");
        end
    endtask

endmodule      counter <= counter + 1'b1;
                end
            end
            else begin
                // Input matches output - reset counter
                counter <= {COUNTER_WIDTH{1'b0}};
            end
        end
    end

endmodule